// Copyright 2015 Heidelberg University Copyright and related rights are
// licensed under the Solderpad Hardware License, Version 0.51 (the "License");
// you may not use this file except in compliance with the License. You may obtain
// a copy of the License at http://solderpad.org/licenses/SHL-0.51. Unless
// required by applicable law or agreed to in writing, software, hardware and
// materials distributed under this License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See
// the License for the specific language governing permissions and limitations
// under the License.


package Sit;
	import Pu_types::*;

	`include "static_mem_model.sv"
	`include "sparse_mem_model.sv"
	`include "state.sv"
	`include "rand_state.sv"
	`include "fixed_state.sv"
	`include "instruction.sv"
	`include "rand_instruction.sv"
	`include "instruction_loader.sv"
	`include "predictor.sv"
	`include "validator.sv"
endpackage
